                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     																								                                                																																																																						                    																																																																																													   																																																																																																																																																																																																																																																																																																																																																																																     																																																																																									                                                                                            																			 													        																																																																																																																																																																																	  			  





  






   

   






																																																																																																																																																																																																																																																																																																																																																																																																																																																						    																																	                        																																																																																																																																																																																																			                      																																																																																																																																																																																																																																																																																																																											    					                                                                                                                                       																																							  													                                                               				                  	           															 																																																																																																														                                                                     																																																																	                                    											             					                                                                                        												  																																															                                                      																																																																																				


   																																																********																																																																																																																																																																				  					                 																																																																																																					       																					  																																			          																		              																																																																																																	           			                                                                                                                                                                                                                                                                                                                                                                                                                                       																													                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     																																									                  	                                        																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																				  																																																																																																																																																																																																																																																																					                      																																																																																																																																																																																																																																																																																																																																																																																																												          													                                                                                   																																																																																																******  																																																		  																																																																			                        																		   																																																																														                                                                                       																																																																																																																																																																																																																																																																																																																																																																																	  																																			******    ****      **    																																																																																																																																																																																				  																										********    ************    																																																					             			             					        		             																																       																																																																																											                                                                                              																				  																														    																																																								  																																			                                                                                    																					                         																																																																																																																														                     										         														                                                                                            ..  ......                                                                                                                                                                                                                                                                                                                                                              ..  ....                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ..................                                         ...................                                                                                                                    ...................................................          ...............................                                                                                         ......................................................................         ...........                          ..........................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    .......                                                                                                                                                                                                                                                                                     ............................................................................................................................................................................                                                                                                                                                         ..................................................                                     ............................................................................................................................................................................................................................ ....... ........   ...................................................................................................................................................................................................                            ..........                                                                                                                        ..........                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      